module CSR (
    input clk, 
    input rst,

    input funct3,
    input funct7,

    input rs1,
    input write_addr,
    input pc,

);
endmodule