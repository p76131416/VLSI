module Decoder (
    
);
    
endmodule